module Add(S, C, A, B);
    input wire [31:0] A, B;
    output wire [31:0] S;
    output wire C;
    wire C3, C7, C11, C15, C19, C23, C27;
    
    addr_4bit FA4_0(S[3:0], C3, A[3:0], B[3:0], 1'b0),
              FA4_1(S[7:4], C7, A[7:4], B[7:4], C3),
              FA4_2(S[11:8], C11, A[11:8], B[11:8], C7),
              FA4_3(S[15:12], C15, A[15:12], B[15:12], C11),
              FA4_4(S[19:16], C19, A[19:16], B[19:16], C15),
              FA4_5(S[23:20], C23, A[23:20], B[23:20], C19),
              FA4_6(S[27:24], C27, A[27:24], B[27:24], C23),
              FA4_7(S[31:28], C, A[31:28], B[31:28], C27);
endmodule
